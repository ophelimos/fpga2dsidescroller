// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mux 

// ============================================================
// File Name: AStep_Mux.v
// Megafunction Name(s):
// 			lpm_mux
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 8.0 Build 231 07/10/2008 SP 1 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2008 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module AStep_Mux (
	data0x,
	data1x,
	data2x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	sel,
	result);

	input	[2:0]  data0x;
	input	[2:0]  data1x;
	input	[2:0]  data2x;
	input	[2:0]  data3x;
	input	[2:0]  data4x;
	input	[2:0]  data5x;
	input	[2:0]  data6x;
	input	[2:0]  data7x;
	input	[2:0]  sel;
	output	[2:0]  result;

	wire [2:0] sub_wire0;
	wire [2:0] sub_wire9 = data7x[2:0];
	wire [2:0] sub_wire8 = data5x[2:0];
	wire [2:0] sub_wire7 = data4x[2:0];
	wire [2:0] sub_wire6 = data3x[2:0];
	wire [2:0] sub_wire5 = data2x[2:0];
	wire [2:0] sub_wire4 = data1x[2:0];
	wire [2:0] sub_wire3 = data0x[2:0];
	wire [2:0] result = sub_wire0[2:0];
	wire [2:0] sub_wire1 = data6x[2:0];
	wire [23:0] sub_wire2 = {sub_wire9, sub_wire1, sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4, sub_wire3};

	lpm_mux	lpm_mux_component (
				.sel (sel),
				.data (sub_wire2),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		lpm_mux_component.lpm_size = 8,
		lpm_mux_component.lpm_type = "LPM_MUX",
		lpm_mux_component.lpm_width = 3,
		lpm_mux_component.lpm_widths = 3;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "8"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "3"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "3"
// Retrieval info: USED_PORT: data0x 0 0 3 0 INPUT NODEFVAL data0x[2..0]
// Retrieval info: USED_PORT: data1x 0 0 3 0 INPUT NODEFVAL data1x[2..0]
// Retrieval info: USED_PORT: data2x 0 0 3 0 INPUT NODEFVAL data2x[2..0]
// Retrieval info: USED_PORT: data3x 0 0 3 0 INPUT NODEFVAL data3x[2..0]
// Retrieval info: USED_PORT: data4x 0 0 3 0 INPUT NODEFVAL data4x[2..0]
// Retrieval info: USED_PORT: data5x 0 0 3 0 INPUT NODEFVAL data5x[2..0]
// Retrieval info: USED_PORT: data6x 0 0 3 0 INPUT NODEFVAL data6x[2..0]
// Retrieval info: USED_PORT: data7x 0 0 3 0 INPUT NODEFVAL data7x[2..0]
// Retrieval info: USED_PORT: result 0 0 3 0 OUTPUT NODEFVAL result[2..0]
// Retrieval info: USED_PORT: sel 0 0 3 0 INPUT NODEFVAL sel[2..0]
// Retrieval info: CONNECT: result 0 0 3 0 @result 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 21 data7x 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 18 data6x 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 15 data5x 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 12 data4x 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 9 data3x 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 6 data2x 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 3 data1x 0 0 3 0
// Retrieval info: CONNECT: @data 0 0 3 0 data0x 0 0 3 0
// Retrieval info: CONNECT: @sel 0 0 3 0 sel 0 0 3 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL AStep_Mux.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL AStep_Mux.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL AStep_Mux.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL AStep_Mux.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL AStep_Mux_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL AStep_Mux_bb.v FALSE
// Retrieval info: LIB_FILE: lpm
